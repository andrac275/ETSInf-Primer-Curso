* F:\Dropbox\Universidad Dropbox\1er Curso\2o Cuatri\TCO\Laboratorio\Pract 6\Apartat1\Apartat2.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 16 19:19:26 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Apartat2.net"
.INC "Apartat2.als"


.probe


.END
