* F:\Dropbox\Universidad Dropbox\1er Curso\2o Cuatri\TCO\Laboratorio\Pract 6\Apartat1\Apartat3Triestado.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 16 19:51:57 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Apartat3Triestado.net"
.INC "Apartat3Triestado.als"


.probe


.END
