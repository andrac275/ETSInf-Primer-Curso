* F:\Dropbox\Universidad Dropbox\1er Curso\2o Cuatri\TCO\Laboratorio\Pract 6\Apartat1\Apartat1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Apr 16 18:00:44 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Apartat1.net"
.INC "Apartat1.als"


.probe


.END
