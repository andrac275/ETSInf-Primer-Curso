* E:\Dropbox\Universidad Dropbox\1er Curso\2o Parcial\TCO\Laboratorio\Pract 2\CircuitoPractica2.sch

* Schematics Version 9.1 - Web Update 1
* Tue Feb 18 17:04:26 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "CircuitoPractica2.net"
.INC "CircuitoPractica2.als"


.probe


.END
