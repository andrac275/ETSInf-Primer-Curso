* W:\TCO\prac4\Circuito_Polarizacion.sch

* Schematics Version 9.1 - Web Update 1
* Tue Mar 03 14:27:46 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Circuito_Polarizacion.net"
.INC "Circuito_Polarizacion.als"


.probe


.END
